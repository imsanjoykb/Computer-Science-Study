module myinv(input a,
		output o);
	assign o = ~a;
endmodule
