module myxor2(input a, b,
		output o);
	assign o = a ^ b;
endmodule 